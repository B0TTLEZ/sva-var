```json
[
    {
        "original_code_slice": ".clk_i               ( clk_i                      ),",
        "mutation_code_slice": ".clk_i               (                            ),"
    },
    {
        "original_code_slice": ".rst_ni              ( rst_ni                     ),",
        "mutation_code_slice": ".rst_ni              (                            ),"
    },
    {
        "original_code_slice": ".req_i               ( req_i                      ),",
        "mutation_code_slice": ".req_i               (                            ),"
    },
    {
        "original_code_slice": ".branch_i            ( prefetch_branch            ),",
        "mutation_code_slice": ".branch_i            (                            ),"
    },
    {
        "original_code_slice": ".addr_i              ( prefetch_addr              ),",
        "mutation_code_slice": ".addr_i              (                            ),"
    },
    {
        "original_code_slice": ".ready_i             ( fetch_ready                ),",
        "mutation_code_slice": ".ready_i             (                            ),"
    },
    {
        "original_code_slice": ".valid_o             ( fetch_valid_raw            ),",
        "mutation_code_slice": ".valid_o             (                            ),"
    },
    {
        "original_code_slice": ".rdata_o             ( fetch_rdata                ),",
        "mutation_code_slice": ".rdata_o             (                            ),"
    },
    {
        "original_code_slice": ".addr_o              ( fetch_addr                 ),",
        "mutation_code_slice": ".addr_o              (                            ),"
    },
    {
        "original_code_slice": ".err_o               ( fetch_err                  ),",
        "mutation_code_slice": ".err_o               (                            ),"
    }
]
```
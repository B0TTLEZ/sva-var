```json
[
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 1; i < N; i++)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i <= N; i++)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; i += 2)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; i--)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = N-1; i >= 0; i--)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N-1; i++)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; i += 0)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; i = i)"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; )"
    },
    {
        "original_code_slice": "for (i = 0; i < N; i++)",
        "mutation_code_slice": "for (i = 0; i < N; i += i)"
    }
]
```
```json
[
    {
        "original_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase",
        "mutation_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase"
    },
    {
        "original_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase",
        "mutation_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n    endcase"
    },
    {
        "original_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase",
        "mutation_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase"
    },
    {
        "original_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase",
        "mutation_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase"
    },
    {
        "original_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase",
        "mutation_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase"
    },
    {
        "original_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase",
        "mutation_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase"
    },
    {
        "original_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase",
        "mutation_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase"
    },
    {
        "original_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase",
        "mutation_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase"
    },
    {
        "original_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_JUMP: fetch_addr_n = branch_target_ex_i;\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase",
        "mutation_code_slice": "unique case (pc_mux_internal)\n      PC_BOOT: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n      PC_EXC:  fetch_addr_n = exc_pc;                       // set PC to exception handler\n      PC_ERET: fetch_addr_n = csr_mepc_i;                   // restore PC when returning from EXC\n      PC_DRET: fetch_addr_n = csr_depc_i;\n      // Without branch predictor will never get pc_mux_internal == PC_BP. We still handle no branch\n      // predictor case here to ensure redundant mux logic isn't synthesised.\n      PC_BP:   fetch_addr_n = BranchPredictor ? predict_branch_pc : { boot_addr_i[31:8], 8'h80 };\n      default: fetch_addr_n = { boot_addr_i[31:8], 8'h80 };\n    endcase"
    },
    {
        "original_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n      default:        exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n    endcase",
        "mutation_code_slice": "unique case (exc_pc_mux_i)\n      EXC_PC_EXC:     exc_pc = { csr_mtvec_i[31:8], 8'h00                };\n      EXC_PC_IRQ:     exc_pc = { csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00 };\n      EXC_PC_DBD:     exc_pc = DmHaltAddr;\n      EXC_PC_DBG_EXC: exc_pc = DmExceptionAddr;\n    endcase"
    }
]
```
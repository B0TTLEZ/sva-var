```json
[
    {
        "original_code_slice" : "if (exc_cause.irq_int) begin\n      // All internal interrupts go to the NMI vector\n      irq_vec = ExcCauseIrqNm.lower_cause;\n    end",
        "mutation_code_slice" : "if (exc_cause.irq_int) begin\n      // All internal interrupts go to the NMI vector\n      // removed else"
    },
    {
        "original_code_slice" : "if (ResetAll) begin : g_instr_rdata_ra\n      always_ff @(posedge clk_i or negedge rst_ni) begin\n        if (!rst_ni) begin\n          instr_rdata_id_o         <= '0;\n          instr_rdata_alu_id_o     <= '0;\n          instr_fetch_err_o        <= '0;\n          instr_fetch_err_plus2_o  <= '0;\n          instr_rdata_c_id_o       <= '0;\n          instr_is_compressed_id_o <= '0;\n          illegal_c_insn_id_o      <= '0;\n          pc_id_o                  <= '0;\n        end else if (if_id_pipe_reg_we) begin\n          instr_rdata_id_o         <= instr_out;\n          instr_rdata_alu_id_o     <= instr_out;\n          instr_fetch_err_o        <= instr_err_out;\n          instr_fetch_err_plus2_o  <= if_instr_err_plus2;\n          instr_rdata_c_id_o       <= if_instr_rdata[15:0];\n          instr_is_compressed_id_o <= instr_is_compressed_out;\n          illegal_c_insn_id_o      <= illegal_c_instr_out;\n          pc_id_o                  <= pc_if_o;\n        end\n      end\n    end",
        "mutation_code_slice" : "if (ResetAll) begin : g_instr_rdata_ra\n      always_ff @(posedge clk_i or negedge rst_ni) begin\n        if (!rst_ni) begin\n          instr_rdata_id_o         <= '0;\n          instr_rdata_alu_id_o     <= '0;\n          instr_fetch_err_o        <= '0;\n          instr_fetch_err_plus2_o  <= '0;\n          instr_rdata_c_id_o       <= '0;\n          instr_is_compressed_id_o <= '0;\n          illegal_c_insn_id_o      <= '0;\n          pc_id_o                  <= '0;\n        end else if (if_id_pipe_reg_we) begin\n          instr_rdata_id_o         <= instr_out;\n          // removed else"
    },
    {
        "original_code_slice" : "if (DummyInstructions) begin : gen_dummy_instr\n    // SEC_CM: CTRL_FLOW.UNPREDICTABLE\n    logic        insert_dummy_instr;\n    logic [31:0] dummy_instr_data;\n\n    ibex_dummy_instr #(\n      .RndCnstLfsrSeed (RndCnstLfsrSeed),\n      .RndCnstLfsrPerm (RndCnstLfsrPerm)\n    ) dummy_instr_i (\n      .clk_i                (clk_i),\n      .rst_ni               (rst_ni),\n      .dummy_instr_en_i     (dummy_instr_en_i),\n      .dummy_instr_mask_i   (dummy_instr_mask_i),\n      .dummy_instr_seed_en_i(dummy_instr_seed_en_i),\n      .dummy_instr_seed_i   (dummy_instr_seed_i),\n      .fetch_valid_i        (fetch_valid),\n      .id_in_ready_i        (id_in_ready_i),\n      .insert_dummy_instr_o (insert_dummy_instr),\n      .dummy_instr_data_o   (dummy_instr_data)\n    );\n\n    // Mux between actual instructions and dummy instructions\n    assign instr_out               = insert_dummy_instr ? dummy_instr_data : instr_decompressed;\n    assign instr_is_compressed_out = insert_dummy_instr ? 1'b0 : instr_is_compressed;\n    assign illegal_c_instr_out     = insert_dummy_instr ? 1'b0 : illegal_c_insn;\n    assign instr_err_out           = insert_dummy_instr ? 1'b0 : if_instr_err;\n\n    // Stall the IF stage if we insert a dummy instruction. The dummy will execute between whatever\n    // is currently in the ID stage and whatever is valid from the prefetch buffer this cycle. The\n    // PC of the dummy instruction will match whatever is next from the prefetch buffer.\n    assign stall_dummy_instr = insert_dummy_instr;\n\n    // Register the dummy instruction indication into the ID stage\n    always_ff @(posedge clk_i or negedge rst_ni) begin\n      if (!rst_ni) begin\n        dummy_instr_id_o <= 1'b0;\n      end else if (if_id_pipe_reg_we) begin\n        dummy_instr_id_o <= insert_dummy_instr;\n      end\n    end\n\n  end else begin : gen_no_dummy_instr",
        "mutation_code_slice" : "if (DummyInstructions) begin : gen_dummy_instr\n    // SEC_CM: CTRL_FLOW.UNPREDICTABLE\n    logic        insert_dummy_instr;\n    logic [31:0] dummy_instr_data;\n\n    ibex_dummy_instr #(\n      .RndCnstLfsrSeed (RndCnstLfsrSeed),\n      .RndCnstLfsrPerm (RndCnstLfsrPerm)\n    ) dummy_instr_i (\n      .clk_i                (clk_i),\n      .rst_ni               (rst_ni),\n      .dummy_instr_en_i     (dummy_instr_en_i),\n      .dummy_instr_mask_i   (dummy_instr_mask_i),\n      .dummy_instr_seed_en_i(dummy_instr_seed_en_i),\n      .dummy_instr_seed_i   (dummy_instr_seed_i),\n      .fetch_valid_i        (fetch_valid),\n      .id_in_ready_i        (id_in_ready_i),\n      .insert_dummy_instr_o (insert_dummy_instr),\n      .dummy_instr_data_o   (dummy_instr_data)\n    );\n\n    // Mux between actual instructions and dummy instructions\n    assign instr_out               = insert_dummy_instr ? dummy_instr_data : instr_decompressed;\n    assign instr_is_compressed_out = insert_dummy_instr ? 1'b0 : instr_is_compressed;\n    assign illegal_c_instr_out     = insert_dummy_instr ? 1'b0 : illegal_c_insn;\n    assign instr_err_out           = insert_dummy_instr ? 1'b0 : if_instr_err;\n\n    // Stall the IF stage if we insert a dummy instruction. The dummy will execute between whatever\n    // is currently in the ID stage and whatever is valid from the prefetch buffer this cycle. The\n    // PC of the dummy instruction will match whatever is next from the prefetch buffer.\n    assign stall_dummy_instr = insert_dummy_instr;\n\n    // Register the dummy instruction indication into the ID stage\n    always_ff @(posedge clk_i or negedge rst_ni) begin\n      if (!rst_ni) begin\n        dummy_instr_id_o <= 1'b0;\n      end else if (if_id_pipe_reg_we) begin\n        dummy_instr_id_o <= insert_dummy_instr;\n      end\n    end\n\n    // removed else"
    },
    {
        "original_code_slice" : "if (ResetAll) begin : g_bp_taken_ra\n      always_ff @(posedge clk_i or negedge rst_ni) begin\n        if (!rst_ni) begin\n          instr_bp_taken_q <= '0;\n        end else if (if_id_pipe_reg_we) begin\n          instr_bp_taken_q <= instr_bp_taken_d;\n        end\n      end\n    end else begin : g_bp_taken_nr",
        "mutation_code_slice" : "if (ResetAll) begin : g_bp_taken_ra\n      always_ff @(posedge clk_i or negedge rst_ni) begin\n        if (!rst_ni) begin\n          instr_bp_taken_q <= '0;\n        end else if (if_id_pipe_reg_we) begin\n          instr_bp_taken_q <= instr_bp_taken_d;\n        end\n      end\n      // removed else"
    },
    {
        "original_code_slice" : "if (ICache) begin : gen_icache\n    // Full I-Cache option\n    ibex_icache #(\n      .ICacheECC       (ICacheECC),\n      .ResetAll        (ResetAll),\n      .BusSizeECC      (BusSizeECC),\n      .TagSizeECC      (TagSizeECC),\n      .LineSizeECC     (LineSizeECC)\n    ) icache_i (\n        .clk_i               ( clk_i                      ),\n        .rst_ni              ( rst_ni                     ),\n\n        .req_i               ( req_i                      ),\n\n        .branch_i            ( prefetch_branch            ),\n        .addr_i              ( prefetch_addr              ),\n\n        .ready_i             ( fetch_ready                ),\n        .valid_o             ( fetch_valid_raw            ),\n        .rdata_o             ( fetch_rdata                ),\n        .addr_o              ( fetch_addr                 ),\n        .err_o               ( fetch_err                  ),\n        .err_plus2_o         ( fetch_err_plus2            ),\n\n        .instr_req_o         ( instr_req_o                ),\n        .instr_addr_o        ( instr_addr_o               ),\n        .instr_gnt_i         ( instr_gnt_i                ),\n        .instr_rvalid_i      ( instr_rvalid_i             ),\n        .instr_rdata_i       ( instr_rdata_i[31:0]        ),\n        .instr_err_i         ( instr_err                  ),\n\n        .ic_tag_req_o        ( ic_tag_req_o               ),\n        .ic_tag_write_o      ( ic_tag_write_o             ),\n        .ic_tag_addr_o       ( ic_tag_addr_o              ),\n        .ic_tag_wdata_o      ( ic_tag_wdata_o             ),\n        .ic_tag_rdata_i      ( ic_tag_rdata_i             ),\n        .ic_data_req_o       ( ic_data_req_o              ),\n        .ic_data_write_o     ( ic_data_write_o            ),\n        .ic_data_addr_o      ( ic_data_addr_o             ),\n        .ic_data_wdata_o     ( ic_data_wdata_o            ),\n        .ic_data_rdata_i     ( ic_data_rdata_i            ),\n        .ic_scr_key_valid_i  ( ic_scr_key_valid_i         ),\n        .ic_scr_key_req_o    ( ic_scr_key_req_o           ),\n\n        .icache_enable_i     ( icache_enable_i            ),\n        .icache_inval_i      ( icache_inval_i             ),\n        .busy_o              ( prefetch_busy              ),\n        .ecc_error_o         ( icache_ecc_error_o         )\n    );\n  end else begin : gen_prefetch_buffer",
        "mutation_code_slice" : "if (ICache) begin : gen_icache\n    // Full I-Cache option\n    ibex_icache #(\n      .ICacheECC       (ICacheECC),\n      .ResetAll        (ResetAll),\n      .BusSizeECC      (BusSizeECC),\n      .TagSizeECC      (TagSizeECC),\n      .LineSizeECC     (LineSizeECC)\n    ) icache_i (\n        .clk_i               ( clk_i                      ),\n        .rst_ni              ( rst_ni                     ),\n\n        .req_i               ( req_i                      ),\n\n        .branch_i            ( prefetch_branch            ),\n        .addr_i              ( prefetch_addr              ),\n\n        .ready_i             ( fetch_ready                ),\n        .valid_o             ( fetch_valid_raw            ),\n        .rdata_o             ( fetch_rdata                ),\n        .addr_o              ( fetch_addr                 ),\n        .err_o               ( fetch_err                  ),\n        .err_plus2_o         ( fetch_err_plus2            ),\n\n        .instr_req_o         ( instr_req_o                ),\n        .instr_addr_o        ( instr_addr_o               ),\n        .instr_gnt_i         ( instr_gnt_i                ),\n        .instr_rvalid_i      ( instr_rvalid_i             ),\n        .instr_rdata_i       ( instr_rdata_i[31:0]        ),\n        .instr_err_i         ( instr_err                  ),\n\n        .ic_tag_req_o        ( ic_tag_req_o               ),\n        .ic_tag_write_o      ( ic_tag_write_o             ),\n        .ic_tag_addr_o       ( ic_tag_addr_o              ),\n        .ic_tag_wdata_o      ( ic_tag_wdata_o             ),\n        .ic_tag_rdata_i      ( ic_tag_rdata_i             ),\n        .ic_data_req_o       ( ic_data_req_o              ),\n        .ic_data_write_o     ( ic_data_write_o            ),\n        .ic_data_addr_o      ( ic_data_addr_o             ),\n        .ic_data_wdata_o     ( ic_data_wdata_o            ),\n        .ic_data_rdata_i     ( ic_data_rdata_i            ),\n        .ic_scr_key_valid_i  ( ic_scr_key_valid_i         ),\n        .ic_scr_key_req_o    ( ic_scr_key_req_o           ),\n\n        .icache_enable_i     ( icache_enable_i            ),\n        .icache_inval_i      ( icache_inval_i             ),\n        .busy_o              ( prefetch_busy              ),\n        .ecc_error_o         ( icache_ecc_error_o         )\n    );\n    // removed else"
    },
    {
        "original_code_slice" : "if (PCIncrCheck) begin : g_secure_pc\n    // SEC_CM: PC.CTRL_FLOW.CONSISTENCY\n    logic [31:0] prev_instr_addr_incr, prev_instr_addr_incr_buf;\n    logic        prev_instr_seq_q, prev_instr_seq_d;\n\n    // Do not check for sequential increase after a branch, jump, exception, interrupt or debug\n    // request, all of which will set branch_req. Also do not check after reset or for dummy\n    // instructions.\n    assign prev_instr_seq_d = (prev_instr_seq_q | instr_new_id_d) &\n        ~branch_req & ~if_instr_err & ~stall_dummy_instr;\n\n    always_ff @(posedge clk_i or negedge rst_ni) begin\n      if (!rst_ni) begin\n        prev_instr_seq_q <= 1'b0;\n      end else begin\n        prev_instr_seq_q <= prev_instr_seq_d;\n      end\n    end\n\n    assign prev_instr_addr_incr = pc_id_o + (instr_is_compressed_id_o ? 32'd2 : 32'd4);\n\n    // Buffer anticipated next PC address to ensure optimiser cannot remove the check.\n    prim_buf #(.Width(32)) u_prev_instr_addr_incr_buf (\n      .in_i (prev_instr_addr_incr),\n      .out_o(prev_instr_addr_incr_buf)\n    );\n\n    // Check that the address equals the previous address +2/+4\n    assign pc_mismatch_alert_o = prev_instr_seq_q & (pc_if_o != prev_instr_addr_incr_buf);\n\n  end else begin : g_no_secure_pc",
        "mutation_code_slice" : "if (PCIncrCheck) begin : g_secure_pc\n    // SEC_CM: PC.CTRL_FLOW.CONSISTENCY\n    logic [31:0] prev_instr_addr_incr, prev_instr_addr_incr_buf;\n    logic        prev_instr_seq_q, prev_instr_seq_d;\n\n    // Do not check for sequential increase after a branch, jump, exception, interrupt or debug\n    // request, all of which will set branch_req. Also do not check after reset or for dummy\n    // instructions.\n    assign prev_instr_seq_d = (prev_instr_seq_q | instr_new_id_d) &\n        ~branch_req & ~if_instr_err & ~stall_dummy_instr;\n\n    always_ff @(posedge clk_i or negedge rst_ni) begin\n      if (!rst_ni) begin\n        prev_instr_seq_q <= 1'b0;\n      end else begin\n        prev_instr_seq_q <= prev_instr_seq_d;\n      end\n    end\n\n    assign prev_instr_addr_incr = pc_id_o + (instr_is_compressed_id_o ? 32'd2 : 32'd4);\n\n    // Buffer anticipated next PC address to ensure optimiser cannot remove the check.\n    prim_buf #(.Width(32)) u_prev_instr_addr_incr_buf (\n      .in_i (prev_instr_addr_incr),\n      .out_o(prev_instr_addr_incr_buf)\n    );\n\n    // Check that the address equals the previous address +2/+4\n    assign pc_mismatch
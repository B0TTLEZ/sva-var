```json
[
    {
        "original_code_slice": "logic              instr_valid_id_d, instr_valid_id_q;",
        "mutation_code_slice": "logic              instr_valid_id_d;"
    },
    {
        "original_code_slice": "logic              instr_new_id_d, instr_new_id_q;",
        "mutation_code_slice": "logic              instr_new_id_d;"
    },
    {
        "original_code_slice": "logic              predict_branch_taken;",
        "mutation_code_slice": "// declaration removed"
    },
    {
        "original_code_slice": "logic [31:0]       predict_branch_pc;",
        "mutation_code_slice": "// declaration removed"
    },
    {
        "original_code_slice": "logic        [4:0] irq_vec;",
        "mutation_code_slice": "// declaration removed"
    },
    {
        "original_code_slice": "logic              instr_skid_bp_taken_q;",
        "mutation_code_slice": "// declaration removed"
    },
    {
        "original_code_slice": "logic              instr_skid_valid_q, instr_skid_valid_d;",
        "mutation_code_slice": "logic              instr_skid_valid_d;"
    },
    {
        "original_code_slice": "logic              instr_bp_taken_q, instr_bp_taken_d;",
        "mutation_code_slice": "logic              instr_bp_taken_d;"
    },
    {
        "original_code_slice": "logic              predict_branch_taken_raw;",
        "mutation_code_slice": "// declaration removed"
    },
    {
        "original_code_slice": "logic [31:0]       prev_instr_addr_incr, prev_instr_addr_incr_buf;",
        "mutation_code_slice": "logic [31:0]       prev_instr_addr_incr_buf;"
    }
]
```